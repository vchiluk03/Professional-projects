package enumtype_i2c;
      typedef enum bit { WRITE, READ } i2c_op_t;
endpackage